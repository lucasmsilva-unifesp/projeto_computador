module ROM
#(parameter DATA_WIDTH=32, parameter ADDR_WIDTH=6)
(
	input [(ADDR_WIDTH-1):0] addr,
	input clk, 
	output reg [(DATA_WIDTH-1):0] q
);

	// Declare the ROM variable
	reg [0:DATA_WIDTH-1] rom[0:2**ADDR_WIDTH-1];
	
	reg primeiroclock = 1;

	// Initialize the ROM with $readmemb.  Put the memory contents
	// in the file single_port_rom_init.txt.  Without this file,
	// this design will not compile.

	// See Verilog LRM 1364-2001 Section 17.2.8 for details on the
	// format of this file, or see the "Using $readmemb and $readmemh"
	// template later in this section.

	always @ (posedge clk)
	begin
		if (primeiroclock) begin 
			$readmemb("fatorial.txt", rom, 0, 2**ADDR_WIDTH-1);
			primeiroclock <= 0;
		end
		
		q <= rom[addr];
	end

endmodule
