module rom
#(
	parameter DATA_WIDTH=32, 
	parameter ADDR_WIDTH=9
)
(
	input [ADDR_WIDTH-1:0] addr,
	input clk, 
	output reg [31:0] q
);

	// Declare the ROM variable
	reg [DATA_WIDTH-1:0] ROM[(2**ADDR_WIDTH)-1:0];
	
	//reg primeiroclock = 1;

	// Initialize the ROM with $readmemb.  Put the memory contents
	// in the file single_port_rom_init.txt.  Without this file,
	// this design will not compile.

	// See Verilog LRM 1364-2001 Section 17.2.8 for details on the
	// format of this file, or see the "Using $readmemb and $readmemh"
	// template later in this section.
	
	
initial begin
	ROM[1] = 32'b000001_111110_000000_00000000000000;
	ROM[2] = 32'b000001_111101_000000_00000000000101;
	ROM[3] = 32'b001100_00000000000000000000011111;
	ROM[4] = 32'b010000_00000000000000000000000000;
	ROM[5] = 32'b010000_00000000000000000000000000;
	ROM[6] = 32'b000100_111111_111110_00000000000001;
	ROM[7] = 32'b000001_001011_111110_00000000000010;
	ROM[8] = 32'b000100_000110_001011_00000000000000;
	ROM[9] = 32'b000001_001100_111110_00000000000011;
	ROM[10] = 32'b000100_000111_001100_00000000000000;
	ROM[11] = 32'b000001_001101_111110_00000000000100;
	ROM[12] = 32'b001111_111111_000000_000000_00_000000;
	ROM[13] = 32'b000001_001111_111110_00000000000010;
	ROM[14] = 32'b000011_010000_001111_00000000000000;
	ROM[15] = 32'b000001_010001_111110_00000000000011;
	ROM[16] = 32'b000011_010010_010001_00000000000000;
	ROM[17] = 32'b000000_010011_010000_010010_00_100000;
	ROM[18] = 32'b000111_010100_010011_000000_00_000000;
	ROM[19] = 32'b000001_010101_111110_00000000000100;
	ROM[20] = 32'b000100_010100_010101_00000000000000;
	ROM[21] = 32'b000001_010110_111110_00000000000100;
	ROM[22] = 32'b000011_010111_010110_00000000000000;
	ROM[23] = 32'b000111_000010_010111_000000_00_000000;
	ROM[24] = 32'b000011_011000_111110_00000000000001;
	ROM[25] = 32'b000111_111111_011000_000000_00_000000;
	ROM[26] = 32'b000010_111101_111101_00000000000101;
	ROM[27] = 32'b000011_011000_111110_00000000000000;
	ROM[28] = 32'b000111_111110_011000_000000_00_000000;
	ROM[29] = 32'b001101_000000_111111_000000_00_000000;
	ROM[30] = 32'b010000_00000000000000000000000000;
	ROM[31] = 32'b010000_000000_000000_000000_00000000;
	ROM[32] = 32'b000100_111111_111110_00000000000001;
	ROM[33] = 32'b000001_011001_111110_00000000000010;
	ROM[34] = 32'b000011_011010_011001_00000000000000;
	ROM[35] = 32'b001110_011010_000000_000000_00_000000;
	ROM[36] = 32'b000111_011011_011010_000000_00_000000;
	ROM[37] = 32'b000001_011100_111110_00000000000010;
	ROM[38] = 32'b000100_011011_011100_00000000000000;
	ROM[39] = 32'b000001_011101_111110_00000000000010;
	ROM[40] = 32'b000011_011110_011101_00000000000000;
	ROM[41] = 32'b000111_000110_011110_000000_00_000000;
	ROM[42] = 32'b001111_011110_000000_000000_00_000000;
	ROM[43] = 32'b000001_011111_111110_00000000000011;
	ROM[44] = 32'b000011_100000_011111_00000000000000;
	ROM[45] = 32'b001110_100000_000000_000000_00_000000;
	ROM[46] = 32'b000111_100001_100000_000000_00_000000;
	ROM[47] = 32'b000001_100010_111110_00000000000011;
	ROM[48] = 32'b000100_100001_100010_00000000000000;
	ROM[49] = 32'b000001_100011_111110_00000000000011;
	ROM[50] = 32'b000011_001011_100011_00000000000000;
	ROM[51] = 32'b000111_000110_001011_000000_00_000000;
	ROM[52] = 32'b001111_001011_000000_000000_00_000000;
	ROM[53] = 32'b000001_001100_111110_00000000000100;
	ROM[54] = 32'b000011_001101_001100_00000000000000;
	ROM[55] = 32'b000001_001110_111110_00000000000010;
	ROM[56] = 32'b000011_001111_001110_00000000000000;
	ROM[57] = 32'b000111_000110_001111_000000_00_000000;
	ROM[58] = 32'b000001_010000_111110_00000000000011;
	ROM[59] = 32'b000011_010001_010000_00000000000000;
	ROM[60] = 32'b000111_000111_010001_000000_00_000000;
	ROM[61] = 32'b000100_111110_111101_00000000000000;
	ROM[62] = 32'b000111_111110_111101_000000_00_000000;
	ROM[63] = 32'b000001_111101_111101_00000000000101;
	ROM[64] = 32'b010010_111111_00000000000000000101;
	ROM[65] = 32'b010000_00000000000000000000000000;
	ROM[66] = 32'b000111_010010_000010_000000_00_000000;
	ROM[67] = 32'b000111_010011_010010_000000_00_000000;
	ROM[68] = 32'b000001_010100_111110_00000000000100;
	ROM[69] = 32'b000100_010011_010100_00000000000000;
	ROM[70] = 32'b000001_010101_111110_00000000000100;
	ROM[71] = 32'b000011_010110_010101_00000000000000;
	ROM[72] = 32'b000111_000110_010110_000000_00_000000;
	ROM[73] = 32'b001111_010110_000000_000000_00_000000;
	ROM[74] = 32'b010001_00000000000000000000000000;
end


	always @ (posedge clk)
	begin
		/*
		if (primeiroclock) begin 
			$readmemb("fatorial.txt", rom, 0, 2**ADDR_WIDTH-1);
			
			primeiroclock <= 0;
		end
		*/
		
		q <= ROM[addr];
	end

endmodule
