module rom
#(
	parameter DATA_WIDTH=32, 
	parameter ADDR_WIDTH=9
)
(
	input [ADDR_WIDTH-1:0] addr,
	input clk, 
	output reg [31:0] q
);

	// Declare the ROM variable
	reg [DATA_WIDTH-1:0] ROM[(2**ADDR_WIDTH)-1:0];
	
	//reg primeiroclock = 1;

	// Initialize the ROM with $readmemb.  Put the memory contents
	// in the file single_port_rom_init.txt.  Without this file,
	// this design will not compile.

	// See Verilog LRM 1364-2001 Section 17.2.8 for details on the
	// format of this file, or see the "Using $readmemb and $readmemh"
	// template later in this section.
	
	
initial begin
ROM[1] = 32'b000001_111110_000000_00000000000000;
ROM[2] = 32'b000001_111101_000000_00000000000100;
ROM[3] = 32'b001100_00000000000000000000101111;
ROM[4] = 32'b010000_00000000000000000000000000;
ROM[5] = 32'b010000_000000_000000_000000_00000000;
ROM[6] = 32'b000100_111111_111110_00000000000001;
ROM[7] = 32'b000001_001011_111110_00000000000010;
ROM[8] = 32'b000100_000110_001011_00000000000000;
ROM[9] = 32'b000001_001100_111110_00000000000011;
ROM[10] = 32'b000100_000111_001100_00000000000000;
ROM[11] = 32'b000011_001101_111110_00000000000011;
ROM[12] = 32'b000001_001110_000000_00000000000000;
ROM[13] = 32'b000000_001111_001101_001110_00_101111;
ROM[14] = 32'b001001_001111_000000_00000000000110;
ROM[15] = 32'b010000_00000000000000000000000000;
ROM[16] = 32'b000011_010000_111110_00000000000010;
ROM[17] = 32'b000111_000010_010000_000000_00_000000;
ROM[19] = 32'b001100_00000000000000000000100111;
ROM[20] = 32'b010000_00000000000000000000000000;
ROM[21] = 32'b010000_000000_000000_000000_00000000;
ROM[22] = 32'b000011_010001_111110_00000000000011;
ROM[23] = 32'b000111_000110_010001_000000_00_000000;
ROM[24] = 32'b000011_010010_111110_00000000000010;
ROM[25] = 32'b000011_010011_111110_00000000000010;
ROM[26] = 32'b000011_010100_111110_00000000000011;
ROM[27] = 32'b000000_010101_010011_010100_00_100011;
ROM[28] = 32'b000011_010110_111110_00000000000011;
ROM[29] = 32'b000000_010111_010101_010110_00_100001;
ROM[30] = 32'b000000_011000_010010_010111_00_100010;
ROM[31] = 32'b000111_000111_011000_000000_00_000000;
ROM[32] = 32'b000100_111110_111101_00000000000000;
ROM[33] = 32'b000111_111110_111101_000000_00_000000;
ROM[34] = 32'b000001_111101_111101_00000000000100;
ROM[35] = 32'b010010_111111_00000000000000000101;
ROM[36] = 32'b010000_00000000000000000000000000;
ROM[37] = 32'b000111_011001_000010_000000_00_000000;
ROM[38] = 32'b000111_000010_011001_000000_00_000000;
ROM[39] = 32'b010000_000000_000000_000000_00000000;
ROM[40] = 32'b000011_011010_111110_00000000000001;
ROM[41] = 32'b000111_111111_011010_000000_00_000000;
ROM[42] = 32'b000010_111101_111101_00000000000100;
ROM[43] = 32'b000011_011011_111110_00000000000000;
ROM[44] = 32'b000111_111110_011011_000000_00_000000;
ROM[45] = 32'b001101_000000_111111_000000_00_000000;
ROM[46] = 32'b010000_00000000000000000000000000;
ROM[47] = 32'b010000_000000_000000_000000_00000000;
ROM[48] = 32'b000100_111111_111110_00000000000001;
ROM[49] = 32'b001110_011100_000000_000000_00_000000;
ROM[50] = 32'b000111_011101_011100_000000_00_000000;
ROM[51] = 32'b000100_011101_111110_00000000000010;
ROM[52] = 32'b001110_011110_000000_000000_00_000000;
ROM[53] = 32'b000111_011111_011110_000000_00_000000;
ROM[54] = 32'b000100_011111_111110_00000000000011;
ROM[55] = 32'b000011_100000_111110_00000000000010;
ROM[56] = 32'b000111_000110_100000_000000_00_000000;
ROM[57] = 32'b000011_100001_111110_00000000000011;
ROM[58] = 32'b000111_000111_100001_000000_00_000000;
ROM[59] = 32'b000100_111110_111101_00000000000000;
ROM[60] = 32'b000111_111110_111101_000000_00_000000;
ROM[61] = 32'b000001_111101_111101_00000000000100;
ROM[62] = 32'b010010_111111_00000000000000000101;
ROM[63] = 32'b010000_00000000000000000000000000;
ROM[64] = 32'b000111_100010_000010_000000_00_000000;
ROM[65] = 32'b000111_000110_100010_000000_00_000000;
ROM[66] = 32'b001111_000110_000000_000000_00_000000;
ROM[67] = 32'b010001_00000000000000000000000000;
end


	always @ (posedge clk)
	begin
		/*
		if (primeiroclock) begin 
			$readmemb("fatorial.txt", rom, 0, 2**ADDR_WIDTH-1);
			
			primeiroclock <= 0;
		end
		*/
		
		q <= ROM[addr];
	end

endmodule
